// module jalr_predictor
// import rv32i_types::*;
